module SimpleFixed2 (
    ports
);
    
endmodule